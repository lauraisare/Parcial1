library verilog;
use verilog.vl_types.all;
entity Contador1_vlg_vec_tst is
end Contador1_vlg_vec_tst;
