library verilog;
use verilog.vl_types.all;
entity Semaforo_salida_vlg_vec_tst is
end Semaforo_salida_vlg_vec_tst;
