library verilog;
use verilog.vl_types.all;
entity FrontSensor_vlg_vec_tst is
end FrontSensor_vlg_vec_tst;
