library verilog;
use verilog.vl_types.all;
entity Controlador_semaforo_vlg_vec_tst is
end Controlador_semaforo_vlg_vec_tst;
