library verilog;
use verilog.vl_types.all;
entity Contador5_vlg_vec_tst is
end Contador5_vlg_vec_tst;
