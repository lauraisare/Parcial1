library verilog;
use verilog.vl_types.all;
entity Contador5_vlg_check_tst is
    port(
        contador_out    : in     vl_logic_vector(6 downto 0);
        sampler_rx      : in     vl_logic
    );
end Contador5_vlg_check_tst;
