library verilog;
use verilog.vl_types.all;
entity PagoPeaje_vlg_vec_tst is
end PagoPeaje_vlg_vec_tst;
